version https://git-lfs.github.com/spec/v1
oid sha256:6517352ef173192e09969f0f08ea6e1b8ec4083881b95823a6d0b1de8daf2742
size 1484
